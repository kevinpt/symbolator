component logo is
  port (
    a,b,c : in bit_vector(1 downto 0);
    x,y : out bit_vector(1 downto 0)
  );
end component;
