component scaled is
  port (
    Clock : in  std_ulogic;
    Reset : in  std_ulogic;
    Din   : in  unsigned;
    Dout  : out unsigned
  );
end component;
